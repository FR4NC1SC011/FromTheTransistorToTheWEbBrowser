module eg1(a,b,sel,clk,en,f);
//Inputs - Outputs
input a,b,sel,clk,en;
output f;
wire f;

// Descripcion de los nodos internos
reg net4,net5;
wire net1,net2,net3;

// Descripcion del dis.





endmodule
